module register_block (
    output reg [31:0] read_data1,
    output reg [31:0] read_data2,
    input [31:0] write_data,
    input [5:0] read_reg1,
    input [5:0] read_reg2,
    input [5:0] write_reg,
    input regWrite
);
    
endmodule