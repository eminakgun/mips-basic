module instruction_block (
    output reg [31:0] instruction,
    input [31:0] pc
);
    
endmodule