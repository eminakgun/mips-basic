
`define ALUop_RTYPE 3'b111
`define ALUop_AND 3'b000
`define ALUop_ADD 3'b101
`define ALUop_SUB 3'b110
`define ALUop_OR  3'b001
`define ALUop_LESS 3'b100