module shift_left_2 (
    output reg [31:0] shifted_address,
    input [31:0] address
);
    
endmodule