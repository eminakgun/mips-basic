module alu (
    output reg [31:0] alu_result,
    output reg zero_bit,
    input [31:0] alu_src1,
    input [31:0] alu_src2,
    input [2:0] alu_ctr);
);
    
endmodule